
module LFSR_Checker (
    input  wire clk                                         , // Señal de reloj
    input  wire i_valid                                     , // Señal de validación del generador LFSR
    input  wire i_soft_reset                                , // Reset sincrónico para registrar el valor de i_seed
    input  wire [7:0] i_LFSR                                , // Valor del LFSR del generador
    input  wire i_rst                                       , // Reset asincrónico
    output reg  o_lock                                        // Señal de salida para indicar si el checker está bloqueado
);

    // Declaración de registros para los contadores

    // Inicialización de los registros
    reg [2:0] valid_counter                                         ;  // Contador para valores válidos (hasta 5)
    reg [2:0] invalid_counter                                       ;  // Contador para valores inválidos (hasta 3)
    reg [7:0] LFSR                                                  ;
    //reg [7:0] aux_LFSR                                            ;
    wire feedback = LFSR[7] ^ (LFSR[6:0]==7'b0000000)               ; 
    reg aux_lock                                                    ;
    

    // Lógica secuencial para los contadores y el estado de bloqueo
    always @(posedge clk or posedge i_rst) begin

        if (i_rst) begin
            // Reset asincrónico: Reinicia todos los contadores y desbloquea
            valid_count   <= 3'b000           ;
            invalid_count <= 2'b00            ;
            o_lock        <= 1'b0             ;
            LFSR          <= 8'b00000001      ;
        end 
        
        else  begin
            // Si i_valid está activo, verifica el valor del LFSR
            if(i_soft_reset) begin
                LFSR <= i_LFSR                  ;
            end 
            
            else if (i_valid) begin
                LFSR[0] <= feedback             ;
                LFSR[1] <= LFSR[0] ^ feedback   ;
                LFSR[2] <= LFSR[1]              ;
                LFSR[3] <= LFSR[2]              ;
                LFSR[4] <= LFSR[3]              ;
                LFSR[5] <= LFSR[4] ^ feedback   ;
                LFSR[6] <= LFSR[5] ^ feedback   ;
                LFSR[7] <= LFSR[6]              ;

                //aux_LFSR <= LFSR              ;

                //if(i_LFSR == aux_LFSR) begin //valid
                if(i_LFSR == LFSR) begin //valid
                    $display(" Valid value detected")                                    ;
                    $display(" input LFSR value: %b", i_LFSR)                            ;
                    $display(" LFSR generated by checker value: %b", LFSR)               ;
                    //$display(" NEXT LFSR value: %b", aux_LFSR)    ;
                    valid_counter = valid_counter + 1               ;
                    invalid_counter <= 0                            ;
                    if(valid_counter>= 5) begin
                        aux_lock <= 1                               ;
                        $display("--------------------")            ;
                        $display("Output LOCK: %b", aux_lock)       ;
                        $display("--------------------")            ;
                        valid_counter <= 0                          ;
                    end
                end

                else if (i_LFSR != LFSR) begin //invalid
                         $display("NOT valid value detected");
                         $display(" input LFSR value: %b", i_LFSR)      ;
                         $display(" LFSR value: %b", LFSR)              ;
                         $display(" NEXT LFSR value: %b", aux_LFSR)     ;
                        invalid_counter = invalid_counter + 1           ;
                        valid_counter <= 0                              ;
                        if(invalid_counter>=3) begin
                            aux_lock=0                                  ;
                            $display("--------------------")            ;
                            $display("Output LOCK: %b", aux_lock)       ;
                            $display("--------------------")            ;
                        end
                end
            end
        end
    end    

assign o_lock = aux_lock                                                ;
  
endmodule
